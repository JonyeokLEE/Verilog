module mx8_32bits(a, b, c, d, e, f, g, h, s2, s1, s0, y);

	input [31:0] a, b, c, d, e, f, g, h;
	input s2, s1, s0; //set input
	
	output [31:0] y; //set output
	
	wire [31:0] w0, w1, w2, w3, w4, w5; //set wire
	
	mx2_32bits mx2_32_0(.d0(a), .d1(b), .s(s0), .y(w0));
	mx2_32bits mx2_32_1(.d0(c), .d1(d), .s(s0),.y(w1));
	mx2_32bits mx2_32_2(.d0(e), .d1(f), .s(s0), .y(w2));
	mx2_32bits mx2_32_3(.d0(g), .d1(h), .s(s0),.y(w3));
	mx2_32bits mx2_32_4(.d0(w0), .d1(w1), .s(s1),.y(w4));
	mx2_32bits mx2_32_5(.d0(w2), .d1(w3), .s(s1),.y(w5));
	mx2_32bits mx2_32_6(.d0(w4), .d1(w5), .s(s2),.y(y)); //connect 7 mx2 module
	
endmodule
